`ifndef AXIS_DEFINES
`define AXIS_DEFINES


`define AXI_DATA_W   32
`define CLOCK_PERIOD 10

`endif // !AXIS_DEFINES