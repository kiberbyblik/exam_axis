`ifndef CLOCK_AGENT_IF
`define CLOCK_AGENT_IF

interface clk_agent_if();

  logic clk;
  
endinterface

`endif //!CLOCK_AGENT_IF
